// Top level module for the policy project
module tb_top;

    import uvm_pkg::*;
    initial begin
        run_test();
    end
endmodule : tb_top
