`ifndef __POLICY_BASE_PKG_SV__
`define __POLICY_BASE_PKG_SV__

package policy_base_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "policy_base.sv"
    `include "policy_list.sv"

endpackage : policy_base_pkg
`endif // __POLICY_BASE_PKG_SV__
